module gpredict_index (
    input [3:0] ghr,
    output [3:0] index
);
    assign index = ghr;
endmodule
